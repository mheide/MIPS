library ieee;
use ieee.std_logic_1164.all;

entity SingleWordReg is
	port (
		clk_i : in std_logic;
		rst_i : in std_logic
	);
end entity SingleWordReg;

architecture behaviour of SingleWordReg is

begin


end architecture;